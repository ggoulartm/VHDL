library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity MatAccControlBlock is
	port(
		-- control inputs
		clock, reset: in std_logic;
		iniciar: in std_logic;
		-- control outputs
		pronto: out std_logic;
		memWrEn: out std_logic;
		-- command outputs
		-- COMPLETE
		-- status intputs
		-- COMPLETE
	);	
end entity;

architecture behav of MatAccControlBlock is
--COMPLETE
begin
--COMPLETE
end;